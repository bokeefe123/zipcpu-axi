module hello_world;
  initial begin
    $display("Hello, Verilator!");
    $finish;
  end
endmodule
